LIBRARY ieee;
USE ieee.std_logic_1164.all;
LIBRARY work;
USE work.all;

ENTITY LAB1a IS
	PORT (
		SW		: IN STD_LOGIC_VECTOR(16 DOWNTO 0);                    
		LEDR	: OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END ENTITY LAB1a;

ARCHITECTURE LAB1a_arch OF LAB1a IS
	COMPONENT MUX21_8B IS
		PORT (
			S		: IN STD_LOGIC;
			X,Y		: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			M		: OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
		);
	END COMPONENT MUX21_8B;
BEGIN
	mux0 : MUX21_8B
	PORT MAP (
		S => SW(16),
		X => SW(7 DOWNTO 0),
		Y => SW(15 DOWNTO 8),
		M => LEDR(7 DOWNTO 0)
	);
END ARCHITECTURE LAB1a_arch;

LIBRARY ieee;
USE ieee.std_logic_1164.all;
LIBRARY work;
USE work.all;

ENTITY MUX21_8B IS 
	PORT (
		S		: IN STD_LOGIC;
		X,Y		: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		M		: OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END ENTITY MUX21_8B;

ARCHITECTURE basic OF  MUX21_8B IS
BEGIN
	MUX21_8B_BEHAVIOR : PROCESS (S,X,Y)
	BEGIN 
		IF (S = '1') THEN M <= Y; ELSE m <= X; END IF;
	END PROCESS MUX21_8B_BEHAVIOR;
END ARCHITECTURE basic;