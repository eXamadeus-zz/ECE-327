LIBRARY ieee;
USE ieee.std_logic_1164.all;
LIBRARY work;
USE work.all;

ENTITY LAB1b IS
	-- PORT (
	-- 	SW		: IN STD_LOGIC_VECTOR(17 DOWNTO 0);                    
	-- 	LEDR	: OUT STD_LOGIC_VECTOR(2 DOWNTO 0)
	-- );

	PORT (
		S : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		U : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		V : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		W : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		X : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		Y : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		M : OUT STD_LOGIC_VECTOR(2 DOWNTO 0)
	);
END ENTITY LAB1b;

ARCHITECTURE LAB1b_arch OF LAB1b IS
	COMPONENT MUX31_5x IS
		PORT (
			S			: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
			U,V,W,X,Y	: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
			M			: OUT STD_LOGIC_VECTOR(2 DOWNTO 0)
		);
	END COMPONENT MUX31_5x;
BEGIN
	mux0 : MUX31_5x
	PORT MAP ( S,U,V,W,X,Y,M
		-- S => SW(17 DOWNTO 15),
		-- U => SW(14 DOWNTO 12),
		-- V => SW(11 DOWNTO 9),
		-- W => SW(8 DOWNTO 6),
		-- X => SW(5 DOWNTO 3),
		-- Y => SW(2 DOWNTO 0),
		-- M => LEDR(2 DOWNTO 0)
	);
END ARCHITECTURE LAB1b_arch;

LIBRARY ieee;
USE ieee.std_logic_1164.all;
LIBRARY work;
USE work.all;

ENTITY MUX31_5x IS 
	PORT (
		S			: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		U,V,W,X,Y	: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		M			: OUT STD_LOGIC_VECTOR(2 DOWNTO 0)
	);
END ENTITY MUX31_5x;

ARCHITECTURE basic OF  MUX31_5x IS
BEGIN
	MUX31_5x_BEHAVIOR : PROCESS (S,U,V,W,X,Y)
	BEGIN 
		CASE S(2 DOWNTO 0) IS
			WHEN "001"  => M <= Y;
			WHEN "010"  => M <= X;
			WHEN "011"  => M <= W;
			WHEN "100"  => M <= V;
			WHEN "101"  => M <= U;
			WHEN OTHERS => M <= "111";
		END CASE;
	END PROCESS MUX31_5x_BEHAVIOR;
END ARCHITECTURE basic;